* Example Testbench Template for IHP SG13G2
* This is a template for creating ngspice testbenches

.title Example Testbench

* Include PDK models
* Update paths according to your PDK installation
.lib '$PDK_ROOT/libs.ref/sg13g2_pr/spice/sg13_lv_models.lib' typical

* Include your design netlist
.include ../schematics/your_block.spice

* Supply voltages
Vdd vdd 0 DC 1.2V
Vss vss 0 DC 0V

* Input stimulus
* Example: Clock signal
Vclk clk 0 PULSE(0 1.2 0 100p 100p 4.9n 10n)

* Example: Reset signal
Vrst rst 0 PULSE(1.2 0 15n 100p 100p 100n 0)

* Example: Enable signal
Ven en 0 PWL(0 0 20n 0 20.1n 1.2 200n 1.2)

* Instantiate your design
X1 clk rst en vdd vss out[0] out[1] out[2] out[3] out[4] out[5] out[6] out[7] carry your_block

* Load capacitance (optional)
.param load_cap=100f
Cout0 out[0] 0 {load_cap}
Cout1 out[1] 0 {load_cap}
Cout2 out[2] 0 {load_cap}
Cout3 out[3] 0 {load_cap}
Cout4 out[4] 0 {load_cap}
Cout5 out[5] 0 {load_cap}
Cout6 out[6] 0 {load_cap}
Cout7 out[7] 0 {load_cap}
Ccarry carry 0 {load_cap}

* Simulation commands
.control
    * Transient analysis
    tran 10p 300n
    
    * Save all signals
    save all
    
    * Plot results
    plot v(clk) v(rst)+2 v(en)+4
    plot v(out[0]) v(out[1])+2 v(out[2])+4 v(out[3])+6
    plot v(out[4]) v(out[5])+2 v(out[6])+4 v(out[7])+6
    plot v(carry)
    
    * Measure propagation delay (example)
    meas tran tpd_rise trig v(clk) val=0.6 rise=10 targ v(out[0]) val=0.6 rise=1
    meas tran tpd_fall trig v(clk) val=0.6 rise=11 targ v(out[0]) val=0.6 fall=1
    
    * Measure power
    meas tran avg_current avg i(Vdd) from=50n to=300n
    let avg_power = avg_current * 1.2
    print avg_power
    
    * Write results
    write example_tb.raw
    
    quit
.endc

.end
